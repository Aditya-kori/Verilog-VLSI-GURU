module h;
initial begin
$display("Hello World");
end
endmodule

//	# Hello World

