module encode(i,y);
input [3:0]i;
output [1:0]y;

