module sample(a,b,c,x,y,z);
	input [7:0]a,b,c;
	output reg[7:0]x,y,z;
	always@(a or b or c) begin
//	x<=a|b;
//	y<=a^b^c;
//	z<=b & ~c;
	x=a|b;
	y=a^b^c;
	z=b & ~c;
	end
endmodule

//# a=21 b=53 c=36 x=53 y=4 z=17
//# a=137 b=94 c=129 x=223 y=86 z=94
//# a=132 b=214 c=9 x=214 y=91 z=214
//# a=240 b=86 c=99 x=246 y=197 z=20
//# a=185 b=123 c=13 x=251 y=207 z=114
//# a=223 b=153 c=141 x=223 y=203 z=16
//# a=194 b=132 c=101 x=198 y=35 z=128
//# a=55 b=82 c=18 x=119 y=119 z=64
//# a=243 b=227 c=1 x=243 y=17 z=226
//# a=215 b=205 c=13 x=223 y=23 z=192


//# a=21 b=53 c=36 x=53 y=4 z=17
//# a=137 b=94 c=129 x=223 y=86 z=94
//# a=132 b=214 c=9 x=214 y=91 z=214
//# a=240 b=86 c=99 x=246 y=197 z=20
//# a=185 b=123 c=13 x=251 y=207 z=114
//# a=223 b=153 c=141 x=223 y=203 z=16
//# a=194 b=132 c=101 x=198 y=35 z=128
//# a=55 b=82 c=18 x=119 y=119 z=64
//# a=243 b=227 c=1 x=243 y=17 z=226
//# a=215 b=205 c=13 x=223 y=23 z=192
