module mux41(s,i,y);
input s[1:0];
input i[3:0];
output y;
assign y=((~s[0])&(~s[1])&i[0])|((s[0])&(~s[1])&i[1])|((~s[0])&(s[1])&i[2])|((s[0])&(s[1])&i[3]);
endmodule


//# s[0]=1 s[1]=0 i0=0 i1=1 i2=0 i3=0 y=1
//# s[0]=0 s[1]=0 i0=0 i1=0 i2=0 i3=1 y=0
//# s[0]=0 s[1]=0 i0=1 i1=0 i2=0 i3=1 y=1
//# s[0]=1 s[1]=0 i0=0 i1=0 i2=1 i3=1 y=0
//# s[0]=0 s[1]=0 i0=1 i1=1 i2=0 i3=1 y=1
//# s[0]=0 s[1]=0 i0=1 i1=1 i2=0 i3=1 y=1
//# s[0]=1 s[1]=0 i0=0 i1=1 i2=0 i3=1 y=1
//# s[0]=0 s[1]=1 i0=0 i1=0 i2=1 i3=0 y=1

