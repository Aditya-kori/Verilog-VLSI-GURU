module mux41(s,i,y);
input s[1:0];
input i[3:0];
reg y0,y1,y2,y3;
output reg y;
always @(*)begin
y0=(~s[0])&(~s[1])&i[0];
y1=(s[0])&(~s[1])&i[1];
y2=(~s[0])&(s[1])&i[2];
y3=(s[0])&(s[1])&i[3];
y=y0|y1|y2|y3;
end
endmodule


//# s[0]=1 s[1]=0 i0=0 i1=1 i2=0 i3=0 y=1
//# s[0]=0 s[1]=0 i0=0 i1=0 i2=0 i3=1 y=0
//# s[0]=0 s[1]=0 i0=1 i1=0 i2=0 i3=1 y=1
//# s[0]=1 s[1]=0 i0=0 i1=0 i2=1 i3=1 y=0
//# s[0]=0 s[1]=0 i0=1 i1=1 i2=0 i3=1 y=1
//# s[0]=0 s[1]=0 i0=1 i1=1 i2=0 i3=1 y=1
//# s[0]=1 s[1]=0 i0=0 i1=1 i2=0 i3=1 y=1
//# s[0]=0 s[1]=1 i0=0 i1=0 i2=1 i3=0 y=1

