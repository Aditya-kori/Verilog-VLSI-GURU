module mux21(s,i0,i1,y);
	input s,i0,i1;
	output y;
endmodule
