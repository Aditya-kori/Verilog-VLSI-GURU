module mux41(s0,s1,i0,i1,i2,i3,y);
input s0,s1,i0,i1,i2,i3;
output y;
assign y=s1?(s0?i3:i2):(s0?i1:i0);
endmodule

//# s1=0,s0=1,i0=0,i1=1,i2=0,i3=0,y=1
//# s1=0,s0=0,i0=0,i1=0,i2=0,i3=1,y=0
//# s1=0,s0=0,i0=1,i1=0,i2=0,i3=1,y=1
//# s1=0,s0=1,i0=0,i1=0,i2=1,i3=1,y=0
//# s1=0,s0=0,i0=1,i1=1,i2=0,i3=1,y=1
//# s1=0,s0=0,i0=1,i1=1,i2=0,i3=1,y=1
//# s1=0,s0=1,i0=0,i1=1,i2=0,i3=1,y=1
//# s1=1,s0=0,i0=0,i1=0,i2=1,i3=0,y=1

